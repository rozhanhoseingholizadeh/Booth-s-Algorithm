`timescale 1ns / 1ps

module Connection_TB;

	// Inputs
	reg CLK;
	reg rx;

	// Outputs
	wire tx;


	reg clken = 1;         // Clock enable signal
   reg [12:0] baud_counter_t = 0; // Baud rate counter
	 
	Connection uut (
		.CLK(CLK), 
		.RX_IN(rx), 
		.TX_OUT(tx)
	);

	initial begin
		CLK = 0;
		rx = 1;

		#70000000;

		// 3 = 0011
		

		//0
		rx = 0;
      #104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;

		#200000;
		
		//0
		rx = 0;
      #104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;

		#200000;

		//1
		rx = 0;
      #104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;

		#200000;


		//1
		rx = 0;
      #104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;

	  #70000000;



		// -7 = 1001

		#200000;

		//1
		rx = 0;
      #104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;

		#200000;
		

		//0
		rx = 0;
      #104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;

		#200000;
		
		//0
		rx = 0;
      #104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;

		#200000;

		//1
		rx = 0;
      #104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 1;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 0;
		#104156.25;
		rx = 1;

		#70000000;
		

	end

	// 50MHz clock
	always @(*)
		#10 CLK <= ~CLK;
		
		
	always @(posedge CLK) begin
		if (baud_counter_t < 2604) begin
			baud_counter_t <= baud_counter_t + 1;
		end else begin
			clken <= ~clken; 
			baud_counter_t <= 0;
		end
	end

	
endmodule

